module wallace(A,B,prod);
input [3:0] A,B;
output [7:0] prod;
   
wire s11,s12,s13,s14,s15,s22,s23,s24,s25,s26,s32,s33,s34,s35,s36,s37;
wire c11,c12,c13,c14,c15,c22,c23,c24,c25,c26,c32,c33,c34,c35,c36,c37;
wire [6:0] p0,p1,p2,p3;

assign  p0 = A & {4{B[0]}};
assign  p1 = A & {4{B[1]}};
assign  p2 = A & {4{B[2]}};
assign  p3 = A & {4{B[3]}};



//first stage
    half_add ha11 (p0[1],p1[0],s11,c11);
    full_add fa12(p0[2],p1[1],p2[0],s12,c12);
    full_add fa13(p0[3],p1[2],p2[1],s13,c13);
    full_add fa14(p1[3],p2[2],p3[1],s14,c14);
    half_add ha15(p2[3],p3[2],s15,c15);

//second stage
    half_add ha22 (c11,s12,s22,c22);
    full_add fa23 (p3[0],c12,s13,s23,c23);
    full_add fa24 (c13,c32,s14,s24,c24);
    full_add fa25 (c14,c24,s15,s25,c25);
    full_add fa26 (c15,c25,p3[3],s26,c26);

//third stage
    half_add ha32(c22,s23,s32,c32);
    half_add ha34(c23,s24,s34,c34);
    half_add ha35(c34,s25,s35,c35);
    half_add ha36(c35,s26,s36,c36);
    half_add ha37(c36,c26,s37,c37);
	 
	 //final product     
assign prod[0] = p0[0];
assign prod[1] = s11;
assign prod[2] = s22;
assign prod[3] = s32;
assign prod[4] = s34;
assign prod[5] = s35;
assign prod[6] = s36;
assign prod[7] = s37;

endmodule